myInstruction_memory_inst : myInstruction_memory PORT MAP (
		address	 => address_sig,
		clock	 => clock_sig,
		q	 => q_sig
	);
